`ifndef DEF_CONFIG
`define DEF_CONFIG

`define RST_PC          64'd0

`endif